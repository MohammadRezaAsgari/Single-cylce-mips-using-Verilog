`timescale 1ns / 1ps

module Add(a, out);
input[7:0] a;
output [7:0] out;

assign out=a+1;

endmodule
